`timescale 1ns/1ns
`include "struct.v"

module struct_tb;
reg a,b,c,d;
wire f,g;

struct uut(a,b,c,d,f,g);
initial begin

	$dumpfile("struct_tb.vcd");
	$dumpvars(0,struct_tb);

	a=0;
	b=0;
	c=0;
	d=0;
	#20;

	a=0;
	b=1;
	c=0;
	d=0;
	#20;

	a=0;
	b=0;
	c=1;
	d=0;
	#20;

	a=0;
	b=0;
	c=0;
	d=1;
	#20;

	a=1;
	b=0;
	c=0;
	d=0;
	#20;


	a=1;
	b=1;
	c=0;
	d=0;
	#20;

	a=1;
	b=0;
	c=1;
	d=0;
	#20;

	a=1;
	b=0;
	c=0;
	d=1;
	#20;

	a=0;
	b=0;
	c=1;
	d=1;
	#20;

	a=0;
	b=1;
	c=0;
	d=1;
	#20;

	a=0;
	b=1;
	c=1;
	d=0;
	#20;


	a=1;
	b=1;
	c=1;
	d=0;
	#20;

	a=1;
	b=1;
	c=0;
	d=1;
	#20;

	a=1;
	b=0;
	c=1;
	d=1;
	#20;

	a=0;
	b=1;
	c=1;
	d=1;
	#20;

	$display("Test Complete");

end


endmodule